`timescale 1ns / 1ps
module seven_seg_decoder(
    input logic [7:0] dataout,
    output logic [6:0] D0, D1, D2, D3, D4, D5, D6, D7
    );

    always_comb
    begin
        D3 = 7'b1111111;
        D4 = 7'b1111111;
        D5 = 7'b1111111;
        D6 = 7'b1111111;
        D7 = 7'b1111111;
        
    case(dataout % 8'd10)   //Ones Digit
        8'd0: D0 = 7'b0000001;//0
        8'd1: D0 = 7'b1001111;//1
        8'd2: D0 = 7'b0010010;//2
        8'd3: D0 = 7'b0000110;//3
        8'd4: D0 = 7'b1001100;//4
        8'd5: D0 = 7'b0100100;//5
        8'd6: D0 = 7'b0100000;//6
        8'd7: D0 = 7'b0001111;//7
        8'd8: D0 = 7'b0000000;//8
        8'd9: D0 = 7'b0000100;//9
        default:D0 = 7'b1111111;
    endcase

    case(dataout /8'd10 % 8'd10)   //tens digit
        8'd0: D1 = 7'b0000001;//0
        8'd1: D1 = 7'b1001111;//1
        8'd2: D1 = 7'b0010010;//2
        8'd3: D1 = 7'b0000110;//3
        8'd4: D1 = 7'b1001100;//4
        8'd5: D1 = 7'b0100100;//5
        8'd6: D1 = 7'b0100000;//6
        8'd7: D1 = 7'b0001111;//7
        8'd8: D1 = 7'b0000000;//8
        8'd9: D1 = 7'b0000100;//9
        default:D1 = 7'b1111111;
    endcase

    case(dataout /8'd100)   //hundreds digit
        8'd0: D2 = 7'b0000001;//0
        8'd1: D2 = 7'b1001111;//1
        8'd2: D2 = 7'b0010010;//2
        8'd3: D2 = 7'b0000110;//3
        8'd4: D2 = 7'b1001100;//4
        8'd5: D2 = 7'b0100100;//5
        8'd6: D2 = 7'b0100000;//6
        8'd7: D2 = 7'b0001111;//7
        8'd8: D2 = 7'b0000000;//8
        8'd9: D2 = 7'b0000100;//9
        default:D2 = 7'b1111111;
    endcase

    end
    
endmodule